--
-- Definition of a single port ROM for KCPSM3 program defined by progctrl.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity progctrl is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end progctrl;
--
architecture low_level_definition of progctrl is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "502E4042502C4045002401540F3E01B601B601B6025601BC01B6C001013D0029";
attribute INIT_01 of ram_1024_x_18  : label is "0F3F01B650F840535003404850E5404950C4404150A54052508E405750494050";
attribute INIT_02 of ram_1024_x_18  : label is "01B60904402F09FEA000C0080006A000016110F0015401424007015401540154";
attribute INIT_03 of ram_1024_x_18  : label is "024F5C3AC902004301540F2E0700080001B6022C01B654414F590154014202F7";
attribute INIT_04 of ram_1024_x_18  : label is "006900594007024F004E020501B6A000011A010D01D0010D0120400703144007";
attribute INIT_05 of ram_1024_x_18  : label is "B0004F0D0142545A4F3A01420E2B404E00796A2B01B60190504E4B04B0004B01";
attribute INIT_06 of ram_1024_x_18  : label is "4B0450744B007BD08D037CD00D2B405D8E01F0E0019712F0014213F0B0004F0A";
attribute INIT_07 of ram_1024_x_18  : label is "C10111A0507920800103010D01E8A00078D0CD0177D0CD01A00079D08D02B400";
attribute INIT_08 of ram_1024_x_18  : label is "01B00321A000011A010D01D05482CA018301A900A8008701010D7130032F010D";
attribute INIT_09 of ram_1024_x_18  : label is "01404007024F01B6009F589801B003311700588E01B01800588E01B01900588E";
attribute INIT_0A of ram_1024_x_18  : label is "01B6170058A501B0180058A501B0190058A501B00321A000011A010D1100010D";
attribute INIT_0B of ram_1024_x_18  : label is "54B8C501018AA900A8008701010301B9051001B9019001B606104007024F00B3";
attribute INIT_0C of ram_1024_x_18  : label is "00D201B6170058A501B0180058A501B0190058A501B00321A00001B654B4C601";
attribute INIT_0D of ram_1024_x_18  : label is "54D8C501018AA900A8008701010301B9051001B9019001B6044606FF4007024F";
attribute INIT_0E of ram_1024_x_18  : label is "0103010D019007000800090001B901540F3D02E901B6A00001B654D4E400C601";
attribute INIT_0F of ram_1024_x_18  : label is "018A010301B6010D01700700080009004007011701B6018A0103070201B9018A";
attribute INIT_10 of ram_1024_x_18  : label is "C720C840C980A000C108400201060106C1080105C720C840C9804007011701B6";
attribute INIT_11 of ram_1024_x_18  : label is "20800103AE008D010D000E00A000010D01FFA000C10801060106C1080100C110";
attribute INIT_12 of ram_1024_x_18  : label is "012A0128A000552BC001000BA00001B6018A10D0018A10E001B6A0000117511C";
attribute INIT_13 of ram_1024_x_18  : label is "C40101380414A0005539C30101330314A0005534C201012E0219A000552FC101";
attribute INIT_14 of ram_1024_x_18  : label is "414C555020084000A000C001514C4F134F014143554720084000C000A000553E";
attribute INIT_15 of ram_1024_x_18  : label is "803AC1015D5BC00A81010130A000CF044154515820014000414C51434F114F01";
attribute INIT_16 of ram_1024_x_18  : label is "02061200B80001677010A000C0F6B80080C6A000A0DFBC00407BB8004061A000";
attribute INIT_17 of ram_1024_x_18  : label is "12000185000E000E000E000E1100A0009200B800016770108101020692000206";
attribute INIT_18 of ram_1024_x_18  : label is "A00001541F1001541F200179A000803A80075988C00AA00011000185A00F1010";
attribute INIT_19 of ram_1024_x_18  : label is "102003060306030603061300B80001A41030A000018A1070018A1080018A1090";
attribute INIT_1A of ram_1024_x_18  : label is "A000800AA000C0F6B80080075DAEC011B800C0E9B80080B9A000D030B80001A4";
attribute INIT_1B of ram_1024_x_18  : label is "01540F5001B601B6A00001540F20A00001540F0DA00001971200002413000024";
attribute INIT_1C of ram_1024_x_18  : label is "01540F6501540F7A01540F6101540F6C01540F4201540F6F01540F6301540F69";
attribute INIT_1D of ram_1024_x_18  : label is "01540F5301540F4101540F4C01540F4601B901540F5201540F4F01540F4E01B9";
attribute INIT_1E of ram_1024_x_18  : label is "0F6D01540F6101540F7201540F6701540F6F01540F7201540F5001B901540F48";
attribute INIT_1F of ram_1024_x_18  : label is "01540F3001540F2E01540F3101540F7601B901540F7201540F6501540F6D0154";
attribute INIT_20 of ram_1024_x_18  : label is "0F6E01540F6901540F7401540F6901540F6101540F57A00001B601B601540F30";
attribute INIT_21 of ram_1024_x_18  : label is "0F5301540F4301540F4D01B901540F7201540F6F01540F6601B901540F670154";
attribute INIT_22 of ram_1024_x_18  : label is "0F6E01540F690243A00001B601540F6501540F6C01540F6901540F4601B90154";
attribute INIT_23 of ram_1024_x_18  : label is "01540F7301540F6501540F7201540F6701540F6F01540F7201540F5001B90154";
attribute INIT_24 of ram_1024_x_18  : label is "01B6A00001B901540F6501540F7301540F6101540F7201540F45A00001B60154";
attribute INIT_25 of ram_1024_x_18  : label is "01540F6C01540F61024301540F2D01540F4501B6A00001B601540F4B01540F4F";
attribute INIT_26 of ram_1024_x_18  : label is "0F6B01540F6301540F6F01540F6C01540F62024301540F2D01540F4201B60154";
attribute INIT_27 of ram_1024_x_18  : label is "0F5001540F2D01540F5001B601540F3301540F2D01540F3101B901540F730154";
attribute INIT_28 of ram_1024_x_18  : label is "01540F57021A01540F6D01540F6101540F7201540F6701540F6F01540F720154";
attribute INIT_29 of ram_1024_x_18  : label is "0F5201B602EE01B901540F6501540F7401540F6901540F7201540F5701540F2D";
attribute INIT_2A of ram_1024_x_18  : label is "01540F3501540F3201B901540F6401540F6101540F6501540F5201540F2D0154";
attribute INIT_2B of ram_1024_x_18  : label is "0F7601540F6501540F4401540F2D01540F4901B601540F7302EE01B901540F36";
attribute INIT_2C of ram_1024_x_18  : label is "01540F4801540F2D01540F4801B602E901B901540F6501540F6301540F690154";
attribute INIT_2D of ram_1024_x_18  : label is "0F6101540F7401540F5301540F2D01540F5301B601540F7001540F6C01540F65";
attribute INIT_2E of ram_1024_x_18  : label is "01540F62A00001540F4401540F49A00001B601540F7301540F7501540F740154";
attribute INIT_2F of ram_1024_x_18  : label is "01540F6601540F6E01540F6F01540F4301B6A00001540F6501540F7401540F79";
attribute INIT_30 of ram_1024_x_18  : label is "01540F6E01540F2F01540F5901540F28024301B901540F6D01540F7201540F69";
attribute INIT_31 of ram_1024_x_18  : label is "01B601540F7401540F7201540F6F01540F6201540F4101B6A00001B901540F29";
attribute INIT_32 of ram_1024_x_18  : label is "01540F3D015401540F7301540F6501540F72015401540F6401540F6101B6A000";
attribute INIT_33 of ram_1024_x_18  : label is "00000000000000000000432E01540F6101540F7401540F6101540F6401B6A000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "43F580016000C004001143FC001353FB20104000E00000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "4DF2118674436CC99F73CFD9FFFEF33FF7C0FF7FCCA2CFFF3DDDDDDDDDF3FFFF";
attribute INITP_01 of ram_1024_x_18 : label is "FF00FFCFF00F3EF5DD5F3F0FF3CF3FBDDD5F3F3FCF3CFEF33FFF3CF3FBCD55C3";
attribute INITP_02 of ram_1024_x_18 : label is "3AA26C668B2662665D4AF4F4F4BD3D3B72DCB72DCB4BCCEF750B2822AA808ABF";
attribute INITP_03 of ram_1024_x_18 : label is "CCCCF3333333333CCCCCF333CCCCCCCCCFB2CB33999D998B2A8B2CCCB3397630";
attribute INITP_04 of ram_1024_x_18 : label is "333CCCF333333CCFCCF33BCCEF33332FCCCCCCCF33BCCCCF333CCCF3333332FC";
attribute INITP_05 of ram_1024_x_18 : label is "CCCCECCCCB32F33333333CCCCCCFF33333333CFCCCF333333FCCCCCCCF333333";
attribute INITP_06 of ram_1024_x_18 : label is "00000000000000000000000000000000003CCCCECF333CCEF33333BCCCCCFCCC";
attribute INITP_07 of ram_1024_x_18 : label is "F233480000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"502E4042502C4045002401540F3E01B601B601B6025601BC01B6C001013D0029",
                INIT_01 => X"0F3F01B650F840535003404850E5404950C4404150A54052508E405750494050",
                INIT_02 => X"01B60904402F09FEA000C0080006A000016110F0015401424007015401540154",
                INIT_03 => X"024F5C3AC902004301540F2E0700080001B6022C01B654414F590154014202F7",
                INIT_04 => X"006900594007024F004E020501B6A000011A010D01D0010D0120400703144007",
                INIT_05 => X"B0004F0D0142545A4F3A01420E2B404E00796A2B01B60190504E4B04B0004B01",
                INIT_06 => X"4B0450744B007BD08D037CD00D2B405D8E01F0E0019712F0014213F0B0004F0A",
                INIT_07 => X"C10111A0507920800103010D01E8A00078D0CD0177D0CD01A00079D08D02B400",
                INIT_08 => X"01B00321A000011A010D01D05482CA018301A900A8008701010D7130032F010D",
                INIT_09 => X"01404007024F01B6009F589801B003311700588E01B01800588E01B01900588E",
                INIT_0A => X"01B6170058A501B0180058A501B0190058A501B00321A000011A010D1100010D",
                INIT_0B => X"54B8C501018AA900A8008701010301B9051001B9019001B606104007024F00B3",
                INIT_0C => X"00D201B6170058A501B0180058A501B0190058A501B00321A00001B654B4C601",
                INIT_0D => X"54D8C501018AA900A8008701010301B9051001B9019001B6044606FF4007024F",
                INIT_0E => X"0103010D019007000800090001B901540F3D02E901B6A00001B654D4E400C601",
                INIT_0F => X"018A010301B6010D01700700080009004007011701B6018A0103070201B9018A",
                INIT_10 => X"C720C840C980A000C108400201060106C1080105C720C840C9804007011701B6",
                INIT_11 => X"20800103AE008D010D000E00A000010D01FFA000C10801060106C1080100C110",
                INIT_12 => X"012A0128A000552BC001000BA00001B6018A10D0018A10E001B6A0000117511C",
                INIT_13 => X"C40101380414A0005539C30101330314A0005534C201012E0219A000552FC101",
                INIT_14 => X"414C555020084000A000C001514C4F134F014143554720084000C000A000553E",
                INIT_15 => X"803AC1015D5BC00A81010130A000CF044154515820014000414C51434F114F01",
                INIT_16 => X"02061200B80001677010A000C0F6B80080C6A000A0DFBC00407BB8004061A000",
                INIT_17 => X"12000185000E000E000E000E1100A0009200B800016770108101020692000206",
                INIT_18 => X"A00001541F1001541F200179A000803A80075988C00AA00011000185A00F1010",
                INIT_19 => X"102003060306030603061300B80001A41030A000018A1070018A1080018A1090",
                INIT_1A => X"A000800AA000C0F6B80080075DAEC011B800C0E9B80080B9A000D030B80001A4",
                INIT_1B => X"01540F5001B601B6A00001540F20A00001540F0DA00001971200002413000024",
                INIT_1C => X"01540F6501540F7A01540F6101540F6C01540F4201540F6F01540F6301540F69",
                INIT_1D => X"01540F5301540F4101540F4C01540F4601B901540F5201540F4F01540F4E01B9",
                INIT_1E => X"0F6D01540F6101540F7201540F6701540F6F01540F7201540F5001B901540F48",
                INIT_1F => X"01540F3001540F2E01540F3101540F7601B901540F7201540F6501540F6D0154",
                INIT_20 => X"0F6E01540F6901540F7401540F6901540F6101540F57A00001B601B601540F30",
                INIT_21 => X"0F5301540F4301540F4D01B901540F7201540F6F01540F6601B901540F670154",
                INIT_22 => X"0F6E01540F690243A00001B601540F6501540F6C01540F6901540F4601B90154",
                INIT_23 => X"01540F7301540F6501540F7201540F6701540F6F01540F7201540F5001B90154",
                INIT_24 => X"01B6A00001B901540F6501540F7301540F6101540F7201540F45A00001B60154",
                INIT_25 => X"01540F6C01540F61024301540F2D01540F4501B6A00001B601540F4B01540F4F",
                INIT_26 => X"0F6B01540F6301540F6F01540F6C01540F62024301540F2D01540F4201B60154",
                INIT_27 => X"0F5001540F2D01540F5001B601540F3301540F2D01540F3101B901540F730154",
                INIT_28 => X"01540F57021A01540F6D01540F6101540F7201540F6701540F6F01540F720154",
                INIT_29 => X"0F5201B602EE01B901540F6501540F7401540F6901540F7201540F5701540F2D",
                INIT_2A => X"01540F3501540F3201B901540F6401540F6101540F6501540F5201540F2D0154",
                INIT_2B => X"0F7601540F6501540F4401540F2D01540F4901B601540F7302EE01B901540F36",
                INIT_2C => X"01540F4801540F2D01540F4801B602E901B901540F6501540F6301540F690154",
                INIT_2D => X"0F6101540F7401540F5301540F2D01540F5301B601540F7001540F6C01540F65",
                INIT_2E => X"01540F62A00001540F4401540F49A00001B601540F7301540F7501540F740154",
                INIT_2F => X"01540F6601540F6E01540F6F01540F4301B6A00001540F6501540F7401540F79",
                INIT_30 => X"01540F6E01540F2F01540F5901540F28024301B901540F6D01540F7201540F69",
                INIT_31 => X"01B601540F7401540F7201540F6F01540F6201540F4101B6A00001B901540F29",
                INIT_32 => X"01540F3D015401540F7301540F6501540F72015401540F6401540F6101B6A000",
                INIT_33 => X"00000000000000000000432E01540F6101540F7401540F6101540F6401B6A000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"43F580016000C004001143FC001353FB20104000E00000000000000000000000",    
               INITP_00 => X"4DF2118674436CC99F73CFD9FFFEF33FF7C0FF7FCCA2CFFF3DDDDDDDDDF3FFFF",
               INITP_01 => X"FF00FFCFF00F3EF5DD5F3F0FF3CF3FBDDD5F3F3FCF3CFEF33FFF3CF3FBCD55C3",
               INITP_02 => X"3AA26C668B2662665D4AF4F4F4BD3D3B72DCB72DCB4BCCEF750B2822AA808ABF",
               INITP_03 => X"CCCCF3333333333CCCCCF333CCCCCCCCCFB2CB33999D998B2A8B2CCCB3397630",
               INITP_04 => X"333CCCF333333CCFCCF33BCCEF33332FCCCCCCCF33BCCCCF333CCCF3333332FC",
               INITP_05 => X"CCCCECCCCB32F33333333CCCCCCFF33333333CFCCCF333333FCCCCCCCF333333",
               INITP_06 => X"00000000000000000000000000000000003CCCCECF333CCEF33333BCCCCCFCCC",
               INITP_07 => X"F233480000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE progctrl.vhd
--
------------------------------------------------------------------------------------
